LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
use IEEE.math_real.all;
ENTITY rom IS
PORT(
	clk : IN std_logic;
	address: IN std_logic_vector(8 DOWNTO 0);
	controlWord: OUT std_logic_vector(25 DOWNTO 0));
END ENTITY rom;

ARCHITECTURE romArch OF rom IS  
	TYPE rom_type IS ARRAY(0 TO 2**9 - 1) of std_logic_vector(25 DOWNTO 0);
	SIGNAL rom : rom_type := (
	--Fetch Instruction
  	0 => "00111011000001100010100001",
  	1 => "01110110000000000001000000",
  	2 => "10001000000000000000000010",
	--Fetch Src Direct
	64 => "00010000010000000000000110",
	--Fetch Src Autoincrement
	72 => "00011011000001100010100101",
	73 => "01110010000000000001000100",
	74 => "10000000010000000000000110",
	--Fetch Src Autodecrement
	80 => "00011010000010100000100101",
	81 => "01110011000000000011000100",
	82 => "10000000010000000000000110",
	--Fectch Src Indexed
	88 => "00111011000001100010100101",
	89 => "01110110000000000000000100",
	90 => "00010000100000000001000100",
	91 => "10001010000001000000000101",
	92 => "01110001000000000010000100",
	93 => "10000000010000000000000110",
	--Fetch Src Direct Indirect
	96 => "00010001000000000011000100",
	97 => "10000000010000000000000110",
	--Fetch Src Autoincrement Indirect
	104 => "00011011000001100010100101",
	105 => "01110010000000000001000100",
	106 => "10000001000000000011000100",
	107 => "10000000010000000000000110",
	--Fetch Src Autodecrement Indirect
	112 => "00011010000010100000100101",
	113 => "01110011000000000011000100",
	114 => "10000001000000000011000100",
	115 => "10000000010000000000000110",
	--Fectch Src Indexed Indirect
	120 => "00111011000001100010100101",
	121 => "01110110000000000000000100",
	122 => "00010000100000000001000100",
	123 => "10001010000001000000000101",
	124 => "01110001000000000010000100",
	125 => "10000001000000000011000100",
	126 => "10000000010000000000000110",
	--Fetch dist Direct
	128 => "00100000100000000000001010",
	--Fetch dist Autoincrement
	136 => "00101011000001100010101001",
	137 => "01110100000000000001001000",
	138 => "10000000100000000000001010",
	--Fetch dist Autodecrement
	144 => "00101010000010100000101001",
	145 => "01110101000000000011001000",
	146 => "10000000100000000000001010",
	--Fetch dist Indexed
	152 => "00111011000001100010101001",
	153 => "01110110000000000000001000",
	154 => "00100000100000000001001000",
	155 => "10001010000001000000001001",
	156 => "01110001000000000010001000",
	157 => "10000000100000000000001010",
	--Fetch dist Direct Indirect
	160 => "00100001000000000011001000",
	161 => "10000000100000000000001010",
	--Fetch dist Autoincrement Indirect
	168 => "00101011000001100010101001",
	169 => "01110100000000000001000100",
	170 => "10000001000000000011001000",
	171 => "10000000100000000000001010",
	--Fetch dist Autodecrement Indirect
	176 => "00101010000010100000101001",
	177 => "01110101000000000011001000",
	178 => "10000001000000000011001000",
	179 => "10000000100000000000001010",
	--Fectch dist Indexed Indirect
	184 => "00111011000001100010101001",
	185 => "01110110000000000000001000",
	186 => "00100000100000000001001000",
	187 => "10001010000001000000001001",
	188 => "01110001000000000010001000",
	189 => "10000001000000000011001000",
	190 => "10000000100000000000001010",
	--ALU Two operand
	192 => "00001010000000100000001110",
	193 => "00001010000001000000001110",
	194 => "00001010000001100000001110",
	195 => "00001010000010000000001110",
	196 => "00001010000010100000001110",
	197 => "00001010000011000000001110",
	198 => "00001010000011100000001110",
	199 => "00001010000100000000001110",
	200 => "00001010000100100000001110",
	--ALU One operand
	256 => "00001010000101000000001110",
	257 => "00001010000101100000001110",
	258 => "00001010000110000000001110",
	259 => "00001010000110100000001110",
	260 => "00001010000111000000001110",
	261 => "00001010000111100000001110",
	262 => "00001010001000000000001110",
	263 => "00001010001000100000001110",
	264 => "00001010001001000000001110",
	--Branch
	320 => "01000000100000000000010000",
	321 => "00111010000001000000010001",
	322 => "01110110000000000000010010",
	--Write
	384 => "01110100000000000000010110",
	385 => "01110000110000000101011010",
	--Zero operand
	448 => "00000000000000001000011110",
	449 => "00000000000000010000011110",
  	OTHERS =>"00000000000000000000000000");
BEGIN
	
        controlWord <= rom(to_integer(unsigned(address)));
    	
END romArch;